***ALU-
.subckt inverter 1 2 3
M1 3 1 2 2 pmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7
.ends

.subckt pass_or 1 2 3 4
M1 2 2 4 4 nmod w=100u l=10u
M2 1 3 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

.subckt pass_and 1 2 3 4
M1 2 3 4 4 nmod w=100u l=10u
M2 1 2 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

.subckt pass_xor 1 2 3 4 5
M1 2 3 5 5 nmod w=100u l=10u
M2 4 1 5 5 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

Va 11 0 dc 0
Vb 12 0 dc 0
Vbin 13 0 dc 0
Vdd 2 0 dc 5V
Xa 11 2 14 inverter
Xb 12 2 15 inverter
Xc 13 2 18 inverter


Xa*b 11 12 14 15 16 pass_xor
X*' 16 2 17 inverter
Xa*b*bin 13 16 17 18 19 pass_xor
Xba' 12 14 11 20 pass_and
Xbin*' 13 17 16 21 pass_and
Xbout 21 20 22 23 pass_or

.tran 0.1m 20m
.control
run
plot V(23)
.endc
.end
