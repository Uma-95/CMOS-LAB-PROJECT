***ALU
.subckt inverter 1 2 3
M1 3 1 2 2 pmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7
.ends

.subckt pass_or 1 2 3 4
M1 2 2 4 4 nmod w=100u l=10u
M2 1 3 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

.subckt pass_and 1 2 3 4
M1 6 5 0 0 nmod w=100u l=10u
M2 6 2 8 8 nmod w=100u l=10u
M3 2 3 4 4 nmod w=100u l=10u
M4 1 2 4 4 nmod w=100u l=10u
M5 2 3 4 4 nmod w=100u l=10u
M6 1 2 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

.subckt pass_xor 1 2 3 4 5
M1 3 1 2 2 pmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7
.ends

Va 11 0 dc 0
Vb 12 0 dc 0
Vc 13 0 dc 0
Vdd 2 0 dc 5V
Xa 11 2 14 inverter
Xb 12 2 15 inverter
Xc 13 2 17 inverter
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7

Xa*b 11 12 14 15 16 pass_xor
Xa*b*c 16 13 18 17 19 pass_xor
X(a*b)c 13 16 18 20 pass_and
Xab 11 12 14 21 pass_and
Xcarry 20 21 22 23 pass_or
M4 24 14 2 2 pmod w=100u l=10u
M5 24 14 0 0 nmod w=100u l=10u
.tran 0.1m 20m
.control
run
plot V(24)
.endc
.end
