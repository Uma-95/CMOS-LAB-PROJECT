***Addition
.subckt inverter 1 2 3
M1 3 1 2 2 pmod w=100u l=10u
M2 3 1 0 0 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7
.ends

.subckt pass_or 1 2 3 4
M1 2 2 4 4 nmod w=100u l=10u
M2 1 3 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends

.subckt pass_and 1 2 3 4
M1 2 3 4 4 nmod w=100u l=10u
M2 1 2 4 4 nmod w=100u l=10u
.model nmod nmos version=54 level=4.7
.ends 

Va 2 0 dc 0
Vb 3 0 dc 0
Vdd 1 0 dc 2V 
Xb 3 1 5 inverter
Xa 2 1 4 inverter
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7
M1 6 5 0 0 nmod w=100u l=10u
M2 8 2 6 6 nmod w=100u l=10u
M3 8 4 7 7 nmod w=100u l=10u
M4 7 3 0 0 nmod w=100u l=10u
M5 8 2 9 9 pmod w=100u l=10u
M6 8 5 9 9 pmod w=100u l=10u
M7 9 4 1 1 pmod w=100u l=10u
M8 9 3 1 1 pmod w=100u l=10u
M9 10 8 1 1 pmod w=100u l=10u
M10 10 8 0 0 nmod w=100u l=10u

.tran 0.1m 20m
.control
run
plot  V(10)
.endc
.end


Vcin 11 0 dc 0
Vdd 1 0 dc 2V 
Xf' 10 1 12 inverter
Xcin' 11 1 13 inverter
.model nmod nmos version=54 level=4.7
.model pmod pmos version=54 level=4.7
M1 14 13 0 0 nmod w=100u l=10u
M2 16 10 14 14 nmod w=100u l=10u
M3 16 12 15 15 nmod w=100u l=10u
M4 15 11 0 0 nmod w=100u l=10u
M5 16 10 17 17 pmod w=100u l=10u
M6 16 13 17 17 pmod w=100u l=10u
M7 17 12 1 1 pmod w=100u l=10u
M8 17 11 1 1 pmod w=100u l=10u
M9 18 16 1 1 pmod w=100u l=10u
M10 18 16 0 0 nmod w=100u l=10u



.tran 0.1m 20m
.control
run
plot  V(18)
.endc
.end
